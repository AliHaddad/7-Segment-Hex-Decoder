module hex_decoder(c, h);
    input [3:0] c;
    output [6:0] h;

    assign h[0] = ~c[3] & ~c[2] & ~c[1] & c[0] |
		~c[3] & c[2] & ~c[1] & ~c[0] |
		c[3] & c[2] & ~c[1] & c[0] |
		c[3] & ~c[2] & c[1] & c[0];

    assign h[1] = c[3] & c[2] & ~c[0] |
		c[3] & c[1] & c[0] |
		c[2] & c[1] & ~c[0] |
		~c[3] & c[2] & ~c[1] & c[0];

    assign h[2] = c[3] & c[2] & ~c[0] |
		c[3] & c[2] & c[1] |
		~c[3] & ~c[2] & c[1] & ~c[0];

    assign h[3] = c[2] & c[1] & c[0] |
		~c[2] & ~c[1] & c[0] |
		~c[3] & c[2] & ~c[1] & ~c[0] |
		c[3] & ~c[2] & c[1] & ~c[0];

    assign h[4] = ~c[3] & c[0] |
		~c[3] & c[2] & ~c[1] |
		~c[2] & ~c[1] & c[0];

    assign h[5] = ~c[3] & ~c[2] & c[0] |
		~c[3] & ~c[2] & c[1] |
		~c[3] & c[1] & c[0] |
		c[3] & c[2] & ~c[1] & c[0];

    assign h[6] = ~c[3] & ~c[2] & ~c[1] |
		~c[3] & c[2] & c[1] & c[0] |
		c[3] & c[2] & ~c[1] & ~c[0];

endmodule
